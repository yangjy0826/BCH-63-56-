//`timescale 1ns / 1ps revised 1
`timescale 1ns / 1ns
module lookuptable(
							     Lookup_Done_1,
							     Lookup_Done_2,
                   clk,
                   rst_n,
                   isEn3,
                   S,
                   s1,
                   s2,
                   p1,
                   p2
//						  p2, revised 9
                   );
  input clk,rst_n,isEn3;
  input [6:0] S;
  input [5:0] s1,s2;
  output [5:0] p1,p2;
  reg [5:0] p1,p2;
  output Lookup_Done_1,Lookup_Done_2;
  reg Lookup_Done_1,Lookup_Done_2;
  
  always@(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
    p1<=6'b0;
    Lookup_Done_1<=1'b0;
    end
    else begin
      if (isEn3==1'b1)  begin
//        if ((!s1)&&(S[0]==1'b1)) begin  /////revised 
//        if ((!s1)&&(s1[0]==1'b1)) begin  /////revised 
        case(s1)
        6'd0:p1<=6'b000000;
        6'd1:p1<=6'b000001;
        6'd2:p1<=6'b000010;
        6'd3:p1<=6'b000111;
        6'd4:p1<=6'b000011;
        6'd5:p1<=6'b001101;
        6'd6:p1<=6'b001000;
        6'd7:p1<=6'b011011;
        6'd8:p1<=6'b000100;
        6'd9:p1<=6'b100001;
        6'd10:p1<=6'b001110;
        6'd11:p1<=6'b100100;
        6'd12:p1<=6'b001001;
        6'd13:p1<=6'b110001;
        6'd14:p1<=6'b011100;
        6'd15:p1<=6'b010011;
        6'd16:p1<=6'b000101;
        6'd17:p1<=6'b011001;
        6'd18:p1<=6'b100010;
        6'd19:p1<=6'b010001;
        6'd20:p1<=6'b001111;
        6'd21:p1<=6'b110101;
        6'd22:p1<=6'b100101;
        6'd23:p1<=6'b110111;
        6'd24:p1<=6'b001010;
        6'd25:p1<=6'b101110;
        6'd26:p1<=6'b110010;
        6'd27:p1<=6'b100111;
        6'd28:p1<=6'b011101;
        6'd29:p1<=6'b101010;
        6'd30:p1<=6'b010100;
        6'd31:p1<=6'b111001;
        6'd32:p1<=6'b000110;
        6'd33:p1<=6'b111111;
        6'd34:p1<=6'b011010;
        6'd35:p1<=6'b001100;
        6'd36:p1<=6'b100011;
        6'd37:p1<=6'b100000;
        6'd38:p1<=6'b010010;
        6'd39:p1<=6'b110000;
        6'd40:p1<=6'b010000;
        6'd41:p1<=6'b011000;
        6'd42:p1<=6'b110110;
        6'd43:p1<=6'b110100;
        6'd44:p1<=6'b100110;
        6'd45:p1<=6'b101101;
        6'd46:p1<=6'b111000;
        6'd47:p1<=6'b101001;
        6'd48:p1<=6'b001011;
        6'd49:p1<=6'b111110;
        6'd50:p1<=6'b101111;
        6'd51:p1<=6'b011111;
        6'd52:p1<=6'b110011;
        6'd53:p1<=6'b010111;
        6'd54:p1<=6'b101000;
        6'd55:p1<=6'b101100;
        6'd56:p1<=6'b011110;
        6'd57:p1<=6'b111101;
        6'd58:p1<=6'b101011;
        6'd59:p1<=6'b010110;
        6'd60:p1<=6'b010101;
        6'd61:p1<=6'b111100;
        6'd62:p1<=6'b111010;
        6'd63:p1<=6'b111011;
        //default: ep<=63'b0;
        endcase  
		  Lookup_Done_1<=1'b1;
      end  
    end
  end
//  end //revised 
  
    always@(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
    p2<=6'b0;
    Lookup_Done_2<=1'b0;
    end
    else begin
      if (isEn3==1'b1) begin
//        if ((!s1)&&(S[0]==1'b1)) begin //// revised 
// if ((!s1)&&(s1[0]==1'b1)) begin  /////revised 
        case(s2)
        6'd0:p2<=6'b000000;
        6'd1:p2<=6'b000001;
        6'd2:p2<=6'b000010;
        6'd3:p2<=6'b000111;
        6'd4:p2<=6'b000011;
        6'd5:p2<=6'b001101;
        6'd6:p2<=6'b001000;
        6'd7:p2<=6'b011011;
        6'd8:p2<=6'b000100;
        6'd9:p2<=6'b100001;
        6'd10:p2<=6'b001110;
        6'd11:p2<=6'b100100;
        6'd12:p2<=6'b001001;
        6'd13:p2<=6'b110001;
        6'd14:p2<=6'b011100;
        6'd15:p2<=6'b010011;
        6'd16:p2<=6'b000101;
        6'd17:p2<=6'b011001;
        6'd18:p2<=6'b100010;
        6'd19:p2<=6'b010001;
        6'd20:p2<=6'b001111;
        6'd21:p2<=6'b110101;
        6'd22:p2<=6'b100101;
        6'd23:p2<=6'b110111;
        6'd24:p2<=6'b001010;
        6'd25:p2<=6'b101110;
        6'd26:p2<=6'b110010;
        6'd27:p2<=6'b100111;
        6'd28:p2<=6'b011101;
        6'd29:p2<=6'b101010;
        6'd30:p2<=6'b010100;
        6'd31:p2<=6'b111001;
        6'd32:p2<=6'b000110;
        6'd33:p2<=6'b111111;
        6'd34:p2<=6'b011010;
        6'd35:p2<=6'b001100;
        6'd36:p2<=6'b100011;
        6'd37:p2<=6'b100000;
        6'd38:p2<=6'b010010;
        6'd39:p2<=6'b110000;
        6'd40:p2<=6'b010000;
        6'd41:p2<=6'b011000;
        6'd42:p2<=6'b110110;
        6'd43:p2<=6'b110100;
        6'd44:p2<=6'b100110;
        6'd45:p2<=6'b101101;
        6'd46:p2<=6'b111000;
        6'd47:p2<=6'b101001;
        6'd48:p2<=6'b001011;
        6'd49:p2<=6'b111110;
        6'd50:p2<=6'b101111;
        6'd51:p2<=6'b011111;
        6'd52:p2<=6'b110011;
        6'd53:p2<=6'b010111;
        6'd54:p2<=6'b101000;
        6'd55:p2<=6'b101100;
        6'd56:p2<=6'b011110;
        6'd57:p2<=6'b111101;
        6'd58:p2<=6'b101011;
        6'd59:p2<=6'b010110;
        6'd60:p2<=6'b010101;
        6'd61:p2<=6'b111100;
        6'd62:p2<=6'b111010;
        6'd63:p2<=6'b111011;
        //default: ep<=63'b0;
        endcase  
		  Lookup_Done_2<=1'b1;
      end  
    end
  end
//  end //evised 
  
endmodule


